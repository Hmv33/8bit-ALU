Time |   A      B     op   | Result  Carry Zero
----------------------------------------------
  10 | 00001010 00000011 000 | 00001101     0     0
  20 | 00001010 00000011 001 | 00000111     0     0
  30 | 00001010 00000011 010 | 00000010     0     0
  40 | 00001010 00000011 011 | 00001011     0     0
  50 | 00001010 00000011 100 | 00001001     0     0
  60 | 00001010 00000000 101 | 11110101     0     0
  70 | 00001010 00000000 110 | 00010100     0     0
  80 | 00001010 00000000 111 | 00000101     0     0
testbench.sv:40: $finish called at 80 (1s)
Done